.MODEL MCERed D
+ IS=5.7909E-12
+ N=3.0457
+ RS=.47801
+ XTI=41.100
+ EG=2.5000

.MODEL MCEGreen D
+ IS=8.5599E-9
+ N=6.9321
+ RS=.61889
+ XTI=62.500
+ EG=2.5000

.MODEL MCEBlue D
+ IS=477.61E-12
+ N=5.7912
+ RS=.56701
+ XTI=62.500
+ EG=2.5000

.MODEL MCEwhite D
+ IS=2.4522E-15
+ N=3.6241
+ RS=.41236
+ XTI=62.500
+ EG=2.5000
